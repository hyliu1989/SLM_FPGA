
module reader_system (
	altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_chipselect,
	altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_address,
	altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_read,
	altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_write,
	altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_byteenable,
	altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_writedata,
	altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_readdata,
	altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_waitrequest,
	altera_up_sd_card_avalon_interface_0_conduit_end_b_SD_cmd,
	altera_up_sd_card_avalon_interface_0_conduit_end_b_SD_dat,
	altera_up_sd_card_avalon_interface_0_conduit_end_b_SD_dat3,
	altera_up_sd_card_avalon_interface_0_conduit_end_o_SD_clock,
	clk_clk,
	sdram_controller_0_wire_addr,
	sdram_controller_0_wire_ba,
	sdram_controller_0_wire_cas_n,
	sdram_controller_0_wire_cke,
	sdram_controller_0_wire_cs_n,
	sdram_controller_0_wire_dq,
	sdram_controller_0_wire_dqm,
	sdram_controller_0_wire_ras_n,
	sdram_controller_0_wire_we_n,
	reset_reset_n,
	sdram_clock_0_clk,
	sdram_controller_0_s1_address,
	sdram_controller_0_s1_byteenable_n,
	sdram_controller_0_s1_chipselect,
	sdram_controller_0_s1_writedata,
	sdram_controller_0_s1_read_n,
	sdram_controller_0_s1_write_n,
	sdram_controller_0_s1_readdata,
	sdram_controller_0_s1_readdatavalid,
	sdram_controller_0_s1_waitrequest);	

	input		altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_chipselect;
	input	[7:0]	altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_address;
	input		altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_read;
	input		altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_write;
	input	[3:0]	altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_byteenable;
	input	[31:0]	altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_writedata;
	output	[31:0]	altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_readdata;
	output		altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_waitrequest;
	inout		altera_up_sd_card_avalon_interface_0_conduit_end_b_SD_cmd;
	inout		altera_up_sd_card_avalon_interface_0_conduit_end_b_SD_dat;
	inout		altera_up_sd_card_avalon_interface_0_conduit_end_b_SD_dat3;
	output		altera_up_sd_card_avalon_interface_0_conduit_end_o_SD_clock;
	input		clk_clk;
	output	[12:0]	sdram_controller_0_wire_addr;
	output	[1:0]	sdram_controller_0_wire_ba;
	output		sdram_controller_0_wire_cas_n;
	output		sdram_controller_0_wire_cke;
	output		sdram_controller_0_wire_cs_n;
	inout	[15:0]	sdram_controller_0_wire_dq;
	output	[1:0]	sdram_controller_0_wire_dqm;
	output		sdram_controller_0_wire_ras_n;
	output		sdram_controller_0_wire_we_n;
	input		reset_reset_n;
	output		sdram_clock_0_clk;
	input	[24:0]	sdram_controller_0_s1_address;
	input	[1:0]	sdram_controller_0_s1_byteenable_n;
	input		sdram_controller_0_s1_chipselect;
	input	[15:0]	sdram_controller_0_s1_writedata;
	input		sdram_controller_0_s1_read_n;
	input		sdram_controller_0_s1_write_n;
	output	[15:0]	sdram_controller_0_s1_readdata;
	output		sdram_controller_0_s1_readdatavalid;
	output		sdram_controller_0_s1_waitrequest;
endmodule
